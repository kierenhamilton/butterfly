module butterfly (
  input Clock, 
  input nReset,           // switch 9
  input [7:0] sswitch,    // switches 0 through 7
  input control,          // switch 8
  );


