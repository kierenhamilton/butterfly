module butterfly_stim; 

timeunit 1ns; 
timeunit 100ps; 

endmodule
